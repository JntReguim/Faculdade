library verilog;
use verilog.vl_types.all;
entity maindec_vlg_vec_tst is
end maindec_vlg_vec_tst;
