library verilog;
use verilog.vl_types.all;
entity aludec_vlg_vec_tst is
end aludec_vlg_vec_tst;
