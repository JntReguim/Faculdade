library verilog;
use verilog.vl_types.all;
entity flopr_vlg_vec_tst is
end flopr_vlg_vec_tst;
