library verilog;
use verilog.vl_types.all;
entity riscvsingle_vlg_vec_tst is
end riscvsingle_vlg_vec_tst;
