library verilog;
use verilog.vl_types.all;
entity dmem_vlg_vec_tst is
end dmem_vlg_vec_tst;
