library verilog;
use verilog.vl_types.all;
entity extend_vlg_vec_tst is
end extend_vlg_vec_tst;
