library verilog;
use verilog.vl_types.all;
entity imem_vlg_vec_tst is
end imem_vlg_vec_tst;
